


 






// file: ibert_7series_gtp_0.v
//////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2012.3
//  \   \         Application : IBERT 7Series 
//  /   /         Filename : example_ibert_7series_gtp_0
// /___/   /\     
// \   \  /  \ 
//  \___\/\___\
//
//
// Module example_ibert_7series_gtp_0
// Generated by Xilinx IBERT_7S 
//////////////////////////////////////////////////////////////////////////////


`define C_NUM_QUADS 1
`define C_REFCLKS_USED 1
module example_ibert_7series_gtp_0
(
  // GT top level ports
  output [(4*`C_NUM_QUADS)-1:0]		TXN_O,
  output [(4*`C_NUM_QUADS)-1:0]		TXP_O,
  input  [(4*`C_NUM_QUADS)-1:0]    	RXN_I,
  input  [(4*`C_NUM_QUADS)-1:0]   	RXP_I,
  input  [`C_REFCLKS_USED-1:0]        	GTREFCLK0P_I,
  input  [`C_REFCLKS_USED-1:0]        	GTREFCLK0N_I,
  input  [`C_REFCLKS_USED-1:0]        	GTREFCLK1P_I,
  input  [`C_REFCLKS_USED-1:0]        	GTREFCLK1N_I,
  output                                txEn,
  input                                 rxLOS,
  input                                 presentb,
  input                                 txFault,
  output  [2:0]                         ledR,
  output  [2:0]                         ledG,
  output  [2:0]                         ledB,
  input                                 jumper8,
  input                                 pllClk,
  input                                 lan9254Clk
);

  //
  // Ibert refclk internal signals
  //
  wire   [`C_NUM_QUADS-1:0]        	gtrefclk0_i;
  wire   [`C_NUM_QUADS-1:0]        	gtrefclk1_i;
  wire   [`C_REFCLKS_USED-1:0]        	refclk0_i;
  wire   [`C_REFCLKS_USED-1:0]        	refclk1_i;
  wire                            	sysclk_i;
  wire                              lanClk_i;
  wire                              pllClk_i;
  
  reg    [24 : 0]                   lanCnt = 0;
  reg    [24 : 0]                   pllCnt = 0;
  reg    [25 : 0]                   refCnt = 0;


  BUFG u_lanclk_bufg( .I( lan9254Clk ), .O (lanClk_i) );
  BUFG u_pllclk_bufg( .I( pllClk     ), .O (pllClk_i) );
  
  always @(posedge lanClk_i) begin
    lanCnt <= lanCnt + 1;
  end
  
  always @(posedge pllClk_i) begin
    pllCnt <= pllCnt + 1;
  end
  
  always @(posedge sysclk_i) begin
    refCnt <= refCnt + 1;
  end
  
  // Refclk IBUFDS instantiations
  //

    IBUFDS_GTE2 u_buf_q0_clk0
      (
        .O            (refclk0_i[0]),
        .ODIV2        (),
        .CEB          (1'b0),
        .I            (GTREFCLK0P_I[0]),
        .IB           (GTREFCLK0N_I[0])
      );

    IBUFDS_GTE2 u_buf_q0_clk1
      (
        .O            (refclk1_i[0]),
        .ODIV2        (),
        .CEB          (1'b0),
        .I            (GTREFCLK1P_I[0]),
        .IB           (GTREFCLK1N_I[0])
      );

  //
  // Refclk connection from each IBUFDS to respective quads depending on the source selected in gui
  //
  assign gtrefclk0_i[0] = refclk0_i[0];
  assign gtrefclk1_i[0] = refclk1_i[0];
  
  assign txEn           = jumper8;
  assign ledB[2]        = presentb;
  assign ledG[2]        = txFault;
  assign ledR[2]        = rxLOS;
  
  assign ledB[1]        = refCnt[25];
  assign ledG[1]        = lanCnt[24];
  assign ledR[1]        = pllCnt[24];
  

  BUFG u_buf_sysclk
    (
      .I              (refclk1_i[0]),
      .O              (sysclk_i)
    );

  //
  // IBERT core instantiation
  //
  ibert_7series_gtp_0 u_ibert_core
    (
      .TXN_O(TXN_O),
      .TXP_O(TXP_O),
      .RXN_I(RXN_I),
      .RXP_I(RXP_I),
      .SYSCLK_I(sysclk_i),
      .GTREFCLK0_I(gtrefclk0_i),
      .GTREFCLK1_I(gtrefclk1_i)
    );

endmodule
